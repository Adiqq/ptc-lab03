library verilog;
use verilog.vl_types.all;
entity licznik7943 is
    port(
        pin_name2       : out    vl_logic;
        pin_name1       : in     vl_logic;
        pin_name3       : out    vl_logic;
        pin_name4       : out    vl_logic;
        pin_name5       : out    vl_logic;
        pin_name6       : out    vl_logic;
        pin_name7       : out    vl_logic;
        pin_name8       : out    vl_logic;
        pin_name9       : out    vl_logic
    );
end licznik7943;
