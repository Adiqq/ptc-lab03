library verilog;
use verilog.vl_types.all;
entity asyncmod12_vlg_vec_tst is
end asyncmod12_vlg_vec_tst;
