library verilog;
use verilog.vl_types.all;
entity licznik74161_vlg_vec_tst is
end licznik74161_vlg_vec_tst;
