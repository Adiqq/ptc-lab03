library verilog;
use verilog.vl_types.all;
entity rewersyjny_vlg_vec_tst is
end rewersyjny_vlg_vec_tst;
