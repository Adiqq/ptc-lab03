library verilog;
use verilog.vl_types.all;
entity rewersyjny_vlg_check_tst is
    port(
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        pin_name7       : in     vl_logic;
        pin_name8       : in     vl_logic;
        pin_name9       : in     vl_logic;
        pin_name10      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end rewersyjny_vlg_check_tst;
