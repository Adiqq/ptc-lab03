library verilog;
use verilog.vl_types.all;
entity licznik7943_vlg_vec_tst is
end licznik7943_vlg_vec_tst;
