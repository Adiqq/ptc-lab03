library verilog;
use verilog.vl_types.all;
entity licznik74163_vlg_vec_tst is
end licznik74163_vlg_vec_tst;
