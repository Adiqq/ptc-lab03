library verilog;
use verilog.vl_types.all;
entity CW4_vlg_vec_tst is
end CW4_vlg_vec_tst;
