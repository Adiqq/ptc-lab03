library verilog;
use verilog.vl_types.all;
entity licznik74193_vlg_vec_tst is
end licznik74193_vlg_vec_tst;
